library verilog;
use verilog.vl_types.all;
entity RV32I_System_tb is
end RV32I_System_tb;
